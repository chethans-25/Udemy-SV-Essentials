/*Generate values between 0 to 7 for addr signal when wr is high and values between 8 to 15 when wr is low. 
Generator code is mentioned in the Instruction tab. 
Verify your code for 20 iterations by sending values of both wr and addr on a console.
*/
